module queue (

input logic data_in,
input logic enqueue_in,
input logic dequeue_in,
input logic reset,
input logic clock_10KHZ,
output logic [7:0] len_out,
output logic [7:0] data_out,

);

logic [7:0] fila [7:0];







endmodule